
module sources_probes (
	source,
	probe,
	source_clk);	

	output	[0:0]	source;
	input	[30:0]	probe;
	input		source_clk;
endmodule
